-- Chris Geraldpaulraj FPGA Final Project 
--- Top Level  Main Entity of whole project.

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.all;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY pr1 IS
	PORT(START: IN STD_LOGIC;
		  RESET: IN STD_LOGIC;
		  CLK: IN STD_LOGIC;
		  VGA_CLK: IN STD_LOGIC;
		  LEFTBUTTON : IN STD_LOGIC;
        RIGHTBUTTON : IN STD_LOGIC;	
		  VGA_HS :   OUT STD_LOGIC;
		  VGA_VS :   OUT STD_LOGIC;
		  VGA_RGB : OUT STD_LOGIC_VECTOR(2 DOWNTO 0)
		 );
		 
END ENTITY;

	ARCHITECTURE RTL OF PR1 IS
	
		COMPONENT ObjAnimation
			PORT(CLK:   IN STD_LOGIC;	
				  HORIZONTAL_CONTROL: IN STD_LOGIC_VECTOR(9 DOWNTO 0);
				  LEFTBUTTON : IN STD_LOGIC;
				  RIGHTBUTTON : IN STD_LOGIC;
				  VERTICAL_CONTROL: IN STD_LOGIC_VECTOR(9 DOWNTO 0);	
				  VIDEO_START : IN STD_LOGIC;
				  VGA_RGB : OUT STD_LOGIC_VECTOR(2 DOWNTO 0)
				 );
				 
		END COMPONENT;
		
		COMPONENT VgaController
			PORT(CLK:   IN STD_LOGIC;
				  RESET: IN STD_LOGIC;	
				  START: IN STD_LOGIC;
				  VERTICAL_CONTROL: OUT STD_LOGIC_VECTOR(9 DOWNTO 0);	
				  HORIZONTAL_CONTROL: OUT STD_LOGIC_VECTOR(9 DOWNTO 0);
				  VGA_HS :   OUT STD_LOGIC;
				  VGA_VS :   OUT STD_LOGIC;
				  VIDEO_START : OUT STD_LOGIC
				  );
				  
		END COMPONENT;
		
		SIGNAL X,Y :  STD_LOGIC_VECTOR(9 DOWNTO 0);
		SIGNAL VIDEO : STD_LOGIC;
		
	BEGIN	
	
		Z_1: ObjAnimation PORT MAP( CLK => CLK , HORIZONTAL_CONTROL => X, LEFTBUTTON => LEFTBUTTON ,RIGHTBUTTON => RIGHTBUTTON, 
                                                         VERTICAL_CONTROL => Y, VIDEO_START => VIDEO , VGA_RGB => VGA_RGB );

		Z_2: VgaController PORT MAP( CLK => CLK, RESET => RESET, START => START, VERTICAL_CONTROL => Y, HORIZONTAL_CONTROL => X ,
                                                             VGA_HS => VGA_HS , VGA_VS => VGA_VS, VIDEO_START => VIDEO );
	
	END RTL;
