--- Creates the animation of the project

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY ObjAnimation IS 
	PORT (CLK : IN STD_LOGIC;
         HORIZONTAL_CONTROL : IN STD_LOGIC_VECTOR(9 DOWNTO 0);
         LEFTBUTTON : IN STD_LOGIC;
         RIGHTBUTTON : IN STD_LOGIC;
         VERTICAL_CONTROL : IN STD_LOGIC_VECTOR(9 DOWNTO 0);
         VIDEO_START : IN STD_LOGIC;
         VGA_RGB : OUT STD_LOGIC_VECTOR(2 DOWNTO 0)
		);
			
END ENTITY;

ARCHITECTURE RTL OF ObjAnimation IS

	TYPE BRICKS IS ARRAY (0 TO 2, 0 TO 9) OF STD_LOGIC;
	SIGNAL BRICKARRAY : BRICKS := ("1111111111", "1111111111", "1111111111");

--- DRAWS THE PADDLE:

	SIGNAL BAR,BAR_NEXT: INTEGER:= 95; --- DISTANCE BETWEEN BAR AND LEFT SIDE OF SCREEN
	CONSTANT BAR_DT: INTEGER:= 400; --- DISTANCE BETWEEN BAR AND TOP SIDE OF SCREEN
	CONSTANT BAR_THICKNESS: INTEGER:= 8; --- THICKNESS OF BAR
	CONSTANT BAR_WIDTH: INTEGER:= 100; --- WIDTH OF BAR
	CONSTANT BAR_SPEED: INTEGER:= 15; --- VELOCITY OF THE BAR
	SIGNAL BAR_START: STD_LOGIC;
	SIGNAL VGA_RGB_BAR: STD_LOGIC_VECTOR(2 DOWNTO 0);

--- DRAWS THE BALL:

	SIGNAL BALL,BALL_NEXT: INTEGER := 80; --- DISTANCE BETWEEN BALL AND LEFT SIDE OF SCREEN
	SIGNAL BALL_TOP,BALL_TOP_NEXT: INTEGER :=80; --- DISTANCE BETWEEN BALL AND TOP SIDE OF SCREEN
	CONSTANT BALL_HEIGHT: INTEGER :=8; --- HEIGHT OF BALL
	CONSTANT BALL_WIDTH: INTEGER :=8; --- WIDTH OF BALL
	CONSTANT HORIZSPEED,VERTSPEED: INTEGER:=2; --- HORIZONTAL AND VERTICAL SPEEDS OF THE BALL 
	SIGNAL BALL_START: STD_LOGIC;
	SIGNAL VGA_RGB_BALL: STD_LOGIC_VECTOR(2 DOWNTO 0);
	
--- MAKES THE MOVEMENT OF PADDLE AND THE BALL:

	SIGNAL RESETREG, RESETREG_NEXT: INTEGER;
	CONSTANT RESET_CONSTANT: INTEGER := 810000;
	SIGNAL RESET_TICK: STD_LOGIC;
	
	--- BALL ANIMATION
	
	SIGNAL H_REG,H_NEXT : INTEGER := 3; -- HORIZONTAL SPEED
	SIGNAL V_REG,V_NEXT : INTEGER := 3; -- VERTICAL SPEED

--- X,Y PIXEL CURSOR

	SIGNAL X,Y : INTEGER RANGE 0 TO 650;

--- MUX

	SIGNAL VDBT:STD_LOGIC_VECTOR(2 DOWNTO 0);

--- BUFFER

	SIGNAL VGA_RGB_REG,VGA_RGB_NEXT : STD_LOGIC_VECTOR(2 DOWNTO 0); 

	BEGIN

		--X,Y PIXEL CURSOR
		X <= CONV_INTEGER(HORIZONTAL_CONTROL);
		Y <= CONV_INTEGER(VERTICAL_CONTROL);

		--RESETING
		
		PROCESS(CLK)
		BEGIN
			  IF CLK'EVENT AND CLK = '1' THEN
					 RESETREG <= RESETREG_NEXT; 
			  END IF;
		END PROCESS;
		
		RESETREG_NEXT <= 0 WHEN RESETREG = RESET_CONSTANT ELSE RESETREG+1;
		
		RESET_TICK <= '1' WHEN RESETREG = 0 ELSE '0';
											
	 	--REGISTER PART
		
		PROCESS(CLK)
		BEGIN
			  IF CLK'EVENT AND CLK='1' THEN
					BALL <= BALL_NEXT;
					BALL_TOP <= BALL_TOP_NEXT;
					H_REG <= H_NEXT;
					V_REG <= V_NEXT;
					BAR <= BAR_NEXT;
				END IF;
		END PROCESS;

		--BAR ANIMATION
		
		PROCESS(BAR,RESET_TICK,RIGHTBUTTON,LEFTBUTTON)
		
		BEGIN
		
			 BAR_NEXT <= BAR;
			 IF RESET_TICK = '1' THEN
				 IF LEFTBUTTON = '1' AND BAR > BAR_SPEED THEN 
					 BAR_NEXT <= BAR - BAR_SPEED;
				 ELSIF RIGHTBUTTON = '1' AND BAR < (639 - BAR_SPEED-BAR_WIDTH) THEN
					  BAR_NEXT <= BAR + BAR_SPEED;
				END IF;
			 END IF;
			 
		END PROCESS;

		--BALL ANIMATION
		PROCESS(RESET_TICK,BALL,BALL_TOP,H_REG,V_REG)
		BEGIN
		
			  BALL_NEXT <= BALL;
			  BALL_NEXT <= BALL_TOP;
			  H_NEXT <= H_REG;
			  V_NEXT <= V_REG;
			  
			  IF RESET_TICK = '1' THEN
			  
				  IF BALL_TOP > 400 AND BALL > (BAR - BALL_WIDTH) AND BALL < (BAR + 120) THEN ---THE BALL HITS  
																																																 
					  V_NEXT<= -VERTSPEED ;
					  
				 ELSIF BALL_TOP < 35 THEN--THE BALL HITS THE WALL
					  V_NEXT<= VERTSPEED;
				 END IF;
				 
				 IF BALL < 8 THEN --THE BALL HITS THE LEFT SIDE OF THE SCREEN
					 H_NEXT <= HORIZSPEED;
					 
				 ELSIF BALL > 600 THEN 
					 H_NEXT<= -HORIZSPEED ; --THE BALL HITS THE RIGHT SIDE OF THE SCREEN
				 END IF; 
				 
				 BALL_NEXT <= BALL + H_REG;
				 BALL_TOP_NEXT <= BALL_TOP + V_REG; 
				 
			 END IF;
		END PROCESS;

		--BAR OBJECT

		BAR_START <= '1' WHEN X > BAR AND X < (BAR+BAR_WIDTH) AND Y> BAR_DT AND Y < (BAR_DT+ BAR_THICKNESS) ELSE '0';
		VGA_RGB_BAR<="010"; --- GREEN

		--BALL OBJECT
		
		BALL_START <= '1' WHEN X > BALL AND X < (BALL+BALL_WIDTH) AND Y> BALL_TOP AND Y < (BALL_TOP+ BALL_HEIGHT) ELSE '0';
		VGA_RGB_BALL <= "100"; --- RED

		--BUFFER
		
		PROCESS(CLK)
		BEGIN
			  IF CLK'EVENT AND CLK='1' THEN
					VGA_RGB_REG <= VGA_RGB_NEXT;
			  END IF;
		END PROCESS;

		--MUX
		
		VDBT <= VIDEO_START & BAR_START & BALL_START; 
		WITH VDBT SELECT
			  VGA_RGB_NEXT <= "101" WHEN "100",--BACKGROUND OF THE SCREEN IS MAGENTA
			  VGA_RGB_BAR WHEN "110",
			  VGA_RGB_BALL WHEN "111",
				"000" WHEN OTHERS;
		
		--OUTPUT
		
		VGA_RGB <= VGA_RGB_REG;

	END RTL;
	
	
